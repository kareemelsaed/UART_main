`include "CONFIG_MACROS_Rx.v"
module UART_Rx
(
    input   wire    [4:0]           prescale,
    input   wire                    RX_IN,
    input   wire                    PAR_EN,
    input   wire                    PAR_TYP,
    input   wire                    CLK,
    input   wire                    RST,
    output  wire     [`WIDTH-1:0]     P_DATA,
    output  wire                     data_valid
);

    /////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////////// Internal Signals ///////////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////
	
wire    [4:0]    edge_count;
wire    [3:0]    bit_count;
        
wire    par_error,
        strt_error,
        stp_error,
        data_samp_enable,
        deser_enable,
        stp_chk_enable,
        strt_chk_enable,
        par_chk_enable,
        counter_enable,
        sampled_bit;
		
	/////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////////// FSM Instantiation //////////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////'

FSM U0_FSM(
    .edge_cnt(edge_count),
    .bit_cnt(bit_count),
    .RX_in(RX_IN),
    .par_en(PAR_EN),
    .par_err(par_error),
    .strt_err(strt_error),
    .stp_err(stp_error),
    .prescale(prescale),
    .clk(CLK),
    .rst(RST),
    .data_samp_en(data_samp_enable),
    .deser_en(deser_enable),
    .data_valid(data_valid),
    .stp_chk_en(stp_chk_enable),
    .strt_chk_en(strt_chk_enable),
    .par_chk_en(par_chk_enable),
    .counter_en(counter_enable)
);

    /////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////// data_sampler Instantiation /////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

data_sampling U0_data_sampling(
    .data_in(RX_IN),
    .prescale(prescale),
    .edge_cnt(edge_count),
    .en_sampler(data_samp_enable),
    .clk(CLK),
    .rst(RST),
    .sampled_bit(sampled_bit)
);

    /////////////////////////////////////////////////////////////////////////////////////////////
    ////////////////////////////// edge_bit_counter Instantiation ///////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////
	
edge_bit_counter U0_edge_bit_counter(
    .prescale(prescale),
    .en_counter(counter_enable),
    .clk(CLK),
    .rst(RST),
    .bit_cnt(bit_count),
    .edge_cnt(edge_count),
    .data_valid(data_valid)
);

    /////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////// deserializer Instantiation /////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

deserializer U0_deserializer(
    .sampled_bit(sampled_bit),
    .data_valid(data_valid),
    .deser_en(deser_enable),
    .clk(CLK),
    .rst(RST),
    .p_data(P_DATA)
);

    /////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////// parity_check Instantiation /////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

parity_check U0_parity_check(
    .sampled_bit(sampled_bit),
    .par_typ(PAR_TYP),
    .clk(CLK),
    .rst(RST),
    .par_check_en(par_chk_enable),
    .par_err(par_error)
);

    /////////////////////////////////////////////////////////////////////////////////////////////
    ///////////////////////////////// strt_check Instantiation //////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

strt_check U0_strt_check(
    .sampled_bit(sampled_bit),
    .strt_check_en(strt_chk_enable),
    .strt_err(strt_error)
);

    /////////////////////////////////////////////////////////////////////////////////////////////
    ////////////////////////////////// stp_check Instantiation //////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

stop_check U0_stop_check(
    .sampled_bit(sampled_bit),
    .stop_check_en(stp_chk_enable),
    .stop_err(stp_error)
);   
endmodule
